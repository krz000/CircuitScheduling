module (clk, rst);

input clk, rst;





endmodule
